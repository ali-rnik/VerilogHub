module adder(input in_A[15:0], output out]15:0]);
	assign out = in_A + 16'd4;
endmodule
