module alu(
