module mips(input clk);

endmodule
